module(aDASCSac

    input a
)



endmodule