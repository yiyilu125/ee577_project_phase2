module(aDASCSac

    input a
)

slkjdqwldjqkwjd

jdlldkqwjldk

ldjasldjl

endmodule