module forward_unit();

endmodule