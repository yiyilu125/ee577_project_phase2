module(

    input a
)



endmodule