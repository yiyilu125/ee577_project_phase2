module(

    input a
)

slkjdqwldjqkwjd

jdlldkqwjldk

ldjasldjl

endmodule