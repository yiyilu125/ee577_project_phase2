module hdu(
    
);

endmodule
